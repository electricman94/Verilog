/*
Author: Ryan Pennell
*/
`ifndef _includes_sv_
`define _includes_sv_
`timescale 1 ns/1 ns

//Debug

//Modules
`include "Module.sv"

`endif
