/*
Author: Ryan Pennell
*/
`ifndef _<Name>_sv_
`define _<Name>_sv_

module <Name> #(
)(
  out,
  in,
  clk,
  reset,
  enable
);

  input wire clk, reset, enable;

  always @ (posedge clk)
  begin

  end
endmodule

`endif
