/*
Author: Ryan Pennell
*/
`ifndef _includes_sv_
`define _includes_sv_
`timescale 1 ns/1 ns

//Debug

//Modules
`include "ALU.sv"
`include "Adder.sv"
`include "Decoder.sv"
`include "Enabler.sv"
`include "InstructionFetch.sv"
`include "Memory.sv"
`include "MemoryAccess.sv"
`include "Mux.sv"
`include "Reg.sv"
`include "Regfile.sv"
`include "SignExtension.sv"
`include "WriteBack.sv"

`endif
